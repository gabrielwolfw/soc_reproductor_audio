// socaudio.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module socaudio (
		input  wire        audio_BCLK,            //          audio.BCLK
		output wire        audio_DACDAT,          //               .DACDAT
		input  wire        audio_DACLRCK,         //               .DACLRCK
		input  wire [3:0]  buttons_export,        //        buttons.export
		input  wire        clk_clk,               //            clk.clk
		input  wire        reset_reset_n,         //          reset.reset_n
		output wire [27:0] seven_segments_export  // seven_segments.export
	);

	wire  [31:0] nios_data_master_readdata;                                 // mm_interconnect_0:NIOS_data_master_readdata -> NIOS:d_readdata
	wire         nios_data_master_waitrequest;                              // mm_interconnect_0:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	wire         nios_data_master_debugaccess;                              // NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_data_master_debugaccess
	wire  [15:0] nios_data_master_address;                                  // NIOS:d_address -> mm_interconnect_0:NIOS_data_master_address
	wire   [3:0] nios_data_master_byteenable;                               // NIOS:d_byteenable -> mm_interconnect_0:NIOS_data_master_byteenable
	wire         nios_data_master_read;                                     // NIOS:d_read -> mm_interconnect_0:NIOS_data_master_read
	wire         nios_data_master_readdatavalid;                            // mm_interconnect_0:NIOS_data_master_readdatavalid -> NIOS:d_readdatavalid
	wire         nios_data_master_write;                                    // NIOS:d_write -> mm_interconnect_0:NIOS_data_master_write
	wire  [31:0] nios_data_master_writedata;                                // NIOS:d_writedata -> mm_interconnect_0:NIOS_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                          // mm_interconnect_0:NIOS_instruction_master_readdata -> NIOS:i_readdata
	wire         nios_instruction_master_waitrequest;                       // mm_interconnect_0:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	wire  [15:0] nios_instruction_master_address;                           // NIOS:i_address -> mm_interconnect_0:NIOS_instruction_master_address
	wire         nios_instruction_master_read;                              // NIOS:i_read -> mm_interconnect_0:NIOS_instruction_master_read
	wire         nios_instruction_master_readdatavalid;                     // mm_interconnect_0:NIOS_instruction_master_readdatavalid -> NIOS:i_readdatavalid
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;     // mm_interconnect_0:AUDIO_avalon_audio_slave_chipselect -> AUDIO:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;       // AUDIO:readdata -> mm_interconnect_0:AUDIO_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;        // mm_interconnect_0:AUDIO_avalon_audio_slave_address -> AUDIO:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;           // mm_interconnect_0:AUDIO_avalon_audio_slave_read -> AUDIO:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;          // mm_interconnect_0:AUDIO_avalon_audio_slave_write -> AUDIO:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;      // mm_interconnect_0:AUDIO_avalon_audio_slave_writedata -> AUDIO:writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;           // NIOS:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;        // NIOS:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;        // mm_interconnect_0:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;            // mm_interconnect_0:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;               // mm_interconnect_0:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;         // mm_interconnect_0:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;              // mm_interconnect_0:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;          // mm_interconnect_0:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                         // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                       // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_seven_segments_s1_chipselect;            // mm_interconnect_0:SEVEN_SEGMENTS_s1_chipselect -> SEVEN_SEGMENTS:chipselect
	wire  [31:0] mm_interconnect_0_seven_segments_s1_readdata;              // SEVEN_SEGMENTS:readdata -> mm_interconnect_0:SEVEN_SEGMENTS_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_segments_s1_address;               // mm_interconnect_0:SEVEN_SEGMENTS_s1_address -> SEVEN_SEGMENTS:address
	wire         mm_interconnect_0_seven_segments_s1_write;                 // mm_interconnect_0:SEVEN_SEGMENTS_s1_write -> SEVEN_SEGMENTS:write_n
	wire  [31:0] mm_interconnect_0_seven_segments_s1_writedata;             // mm_interconnect_0:SEVEN_SEGMENTS_s1_writedata -> SEVEN_SEGMENTS:writedata
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                     // BUTTONS:readdata -> mm_interconnect_0:BUTTONS_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                      // mm_interconnect_0:BUTTONS_s1_address -> BUTTONS:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         irq_mapper_receiver0_irq;                                  // AUDIO:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // TIMER:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios_irq_irq;                                              // irq_mapper:sender_irq -> NIOS:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [AUDIO:reset, BUTTONS:reset_n, JTAG_UART:rst_n, NIOS:reset_n, RAM:reset, SEVEN_SEGMENTS:reset_n, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [NIOS:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	socaudio_AUDIO audio (
		.clk         (clk_clk),                                               //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                              //          interrupt.irq
		.AUD_BCLK    (audio_BCLK),                                            // external_interface.export
		.AUD_DACDAT  (audio_DACDAT),                                          //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                          //                   .export
	);

	socaudio_AUDIO_CLOCK audio_clock (
		.ref_clk_clk        (clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n), //    ref_reset.reset
		.audio_clk_clk      (),               //    audio_clk.clk
		.reset_source_reset ()                // reset_source.reset
	);

	socaudio_BUTTONS buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_export)                         // external_connection.export
	);

	socaudio_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	socaudio_NIOS nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	socaudio_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	socaudio_SEVEN_SEGMENTS seven_segments (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_seven_segments_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_segments_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_segments_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_segments_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_segments_s1_readdata),   //                    .readdata
		.out_port   (seven_segments_export)                           // external_connection.export
	);

	socaudio_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	socaudio_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                             (clk_clk),                                                   //                          CLK_clk.clk
		.NIOS_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                            // NIOS_reset_reset_bridge_in_reset.reset
		.NIOS_data_master_address                (nios_data_master_address),                                  //                 NIOS_data_master.address
		.NIOS_data_master_waitrequest            (nios_data_master_waitrequest),                              //                                 .waitrequest
		.NIOS_data_master_byteenable             (nios_data_master_byteenable),                               //                                 .byteenable
		.NIOS_data_master_read                   (nios_data_master_read),                                     //                                 .read
		.NIOS_data_master_readdata               (nios_data_master_readdata),                                 //                                 .readdata
		.NIOS_data_master_readdatavalid          (nios_data_master_readdatavalid),                            //                                 .readdatavalid
		.NIOS_data_master_write                  (nios_data_master_write),                                    //                                 .write
		.NIOS_data_master_writedata              (nios_data_master_writedata),                                //                                 .writedata
		.NIOS_data_master_debugaccess            (nios_data_master_debugaccess),                              //                                 .debugaccess
		.NIOS_instruction_master_address         (nios_instruction_master_address),                           //          NIOS_instruction_master.address
		.NIOS_instruction_master_waitrequest     (nios_instruction_master_waitrequest),                       //                                 .waitrequest
		.NIOS_instruction_master_read            (nios_instruction_master_read),                              //                                 .read
		.NIOS_instruction_master_readdata        (nios_instruction_master_readdata),                          //                                 .readdata
		.NIOS_instruction_master_readdatavalid   (nios_instruction_master_readdatavalid),                     //                                 .readdatavalid
		.AUDIO_avalon_audio_slave_address        (mm_interconnect_0_audio_avalon_audio_slave_address),        //         AUDIO_avalon_audio_slave.address
		.AUDIO_avalon_audio_slave_write          (mm_interconnect_0_audio_avalon_audio_slave_write),          //                                 .write
		.AUDIO_avalon_audio_slave_read           (mm_interconnect_0_audio_avalon_audio_slave_read),           //                                 .read
		.AUDIO_avalon_audio_slave_readdata       (mm_interconnect_0_audio_avalon_audio_slave_readdata),       //                                 .readdata
		.AUDIO_avalon_audio_slave_writedata      (mm_interconnect_0_audio_avalon_audio_slave_writedata),      //                                 .writedata
		.AUDIO_avalon_audio_slave_chipselect     (mm_interconnect_0_audio_avalon_audio_slave_chipselect),     //                                 .chipselect
		.BUTTONS_s1_address                      (mm_interconnect_0_buttons_s1_address),                      //                       BUTTONS_s1.address
		.BUTTONS_s1_readdata                     (mm_interconnect_0_buttons_s1_readdata),                     //                                 .readdata
		.JTAG_UART_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //      JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                 .write
		.JTAG_UART_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                 .read
		.JTAG_UART_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                 .readdata
		.JTAG_UART_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                 .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.NIOS_debug_mem_slave_address            (mm_interconnect_0_nios_debug_mem_slave_address),            //             NIOS_debug_mem_slave.address
		.NIOS_debug_mem_slave_write              (mm_interconnect_0_nios_debug_mem_slave_write),              //                                 .write
		.NIOS_debug_mem_slave_read               (mm_interconnect_0_nios_debug_mem_slave_read),               //                                 .read
		.NIOS_debug_mem_slave_readdata           (mm_interconnect_0_nios_debug_mem_slave_readdata),           //                                 .readdata
		.NIOS_debug_mem_slave_writedata          (mm_interconnect_0_nios_debug_mem_slave_writedata),          //                                 .writedata
		.NIOS_debug_mem_slave_byteenable         (mm_interconnect_0_nios_debug_mem_slave_byteenable),         //                                 .byteenable
		.NIOS_debug_mem_slave_waitrequest        (mm_interconnect_0_nios_debug_mem_slave_waitrequest),        //                                 .waitrequest
		.NIOS_debug_mem_slave_debugaccess        (mm_interconnect_0_nios_debug_mem_slave_debugaccess),        //                                 .debugaccess
		.RAM_s1_address                          (mm_interconnect_0_ram_s1_address),                          //                           RAM_s1.address
		.RAM_s1_write                            (mm_interconnect_0_ram_s1_write),                            //                                 .write
		.RAM_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                         //                                 .readdata
		.RAM_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                        //                                 .writedata
		.RAM_s1_byteenable                       (mm_interconnect_0_ram_s1_byteenable),                       //                                 .byteenable
		.RAM_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                       //                                 .chipselect
		.RAM_s1_clken                            (mm_interconnect_0_ram_s1_clken),                            //                                 .clken
		.SEVEN_SEGMENTS_s1_address               (mm_interconnect_0_seven_segments_s1_address),               //                SEVEN_SEGMENTS_s1.address
		.SEVEN_SEGMENTS_s1_write                 (mm_interconnect_0_seven_segments_s1_write),                 //                                 .write
		.SEVEN_SEGMENTS_s1_readdata              (mm_interconnect_0_seven_segments_s1_readdata),              //                                 .readdata
		.SEVEN_SEGMENTS_s1_writedata             (mm_interconnect_0_seven_segments_s1_writedata),             //                                 .writedata
		.SEVEN_SEGMENTS_s1_chipselect            (mm_interconnect_0_seven_segments_s1_chipselect),            //                                 .chipselect
		.TIMER_s1_address                        (mm_interconnect_0_timer_s1_address),                        //                         TIMER_s1.address
		.TIMER_s1_write                          (mm_interconnect_0_timer_s1_write),                          //                                 .write
		.TIMER_s1_readdata                       (mm_interconnect_0_timer_s1_readdata),                       //                                 .readdata
		.TIMER_s1_writedata                      (mm_interconnect_0_timer_s1_writedata),                      //                                 .writedata
		.TIMER_s1_chipselect                     (mm_interconnect_0_timer_s1_chipselect)                      //                                 .chipselect
	);

	socaudio_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
